class adder_config extends uvm_object;
	`uvm_object_utils(adder_config);

	function new (string name = "");
		super.new(name);
	endfunction

endclass
