	import uvm_pkg::*;
package adder_package;
	`include "adder_transaction_item.sv"
	`include "adder_sequences.sv"
	`include "adder_driver.sv"
	`include "adder_monitor.sv"
	`include "adder_agent.sv"
	`include "adder_scoreboard.sv"
	`include "adder_env.sv"
	`include "adder_test.sv"
	`include "adder_config.sv"

endpackage
